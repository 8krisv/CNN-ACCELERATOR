// nios_system.v

// Generated using ACDS version 20.1 711

`timescale 1 ps / 1 ps
module nios_system (
		input  wire  clk_clk,                                              //                                      clk.clk
		output wire  cnn_accelerator_avalon_0_control_signals_finished,    // cnn_accelerator_avalon_0_control_signals.finished
		input  wire  cnn_accelerator_avalon_0_control_signals_finished_ok, //                                         .finished_ok
		input  wire  cnn_accelerator_avalon_0_control_signals_same_w,      //                                         .same_w
		input  wire  cnn_accelerator_avalon_0_control_signals_start,       //                                         .start
		input  wire  reset_reset_n                                         //                                    reset.reset_n
	);

	wire  [31:0] cnn_accelerator_avalon_0_avalon_master_readdata;                      // mm_interconnect_0:cnn_accelerator_avalon_0_avalon_master_readdata -> cnn_accelerator_avalon_0:AVS_m0_readdata
	wire         cnn_accelerator_avalon_0_avalon_master_waitrequest;                   // mm_interconnect_0:cnn_accelerator_avalon_0_avalon_master_waitrequest -> cnn_accelerator_avalon_0:AVS_m0_waitrequest
	wire  [17:0] cnn_accelerator_avalon_0_avalon_master_address;                       // cnn_accelerator_avalon_0:AVS_m0_adress -> mm_interconnect_0:cnn_accelerator_avalon_0_avalon_master_address
	wire   [3:0] cnn_accelerator_avalon_0_avalon_master_byteenable;                    // cnn_accelerator_avalon_0:AVS_m0_byteenable -> mm_interconnect_0:cnn_accelerator_avalon_0_avalon_master_byteenable
	wire         cnn_accelerator_avalon_0_avalon_master_read;                          // cnn_accelerator_avalon_0:AVS_m0_read -> mm_interconnect_0:cnn_accelerator_avalon_0_avalon_master_read
	wire         cnn_accelerator_avalon_0_avalon_master_write;                         // cnn_accelerator_avalon_0:AVS_m0_write -> mm_interconnect_0:cnn_accelerator_avalon_0_avalon_master_write
	wire  [31:0] cnn_accelerator_avalon_0_avalon_master_writedata;                     // cnn_accelerator_avalon_0:AVS_m0_writedata -> mm_interconnect_0:cnn_accelerator_avalon_0_avalon_master_writedata
	wire         mm_interconnect_0_onchip_d_memory_s2_chipselect;                      // mm_interconnect_0:onchip_d_memory_s2_chipselect -> onchip_d_memory:chipselect2
	wire  [31:0] mm_interconnect_0_onchip_d_memory_s2_readdata;                        // onchip_d_memory:readdata2 -> mm_interconnect_0:onchip_d_memory_s2_readdata
	wire   [9:0] mm_interconnect_0_onchip_d_memory_s2_address;                         // mm_interconnect_0:onchip_d_memory_s2_address -> onchip_d_memory:address2
	wire   [3:0] mm_interconnect_0_onchip_d_memory_s2_byteenable;                      // mm_interconnect_0:onchip_d_memory_s2_byteenable -> onchip_d_memory:byteenable2
	wire         mm_interconnect_0_onchip_d_memory_s2_write;                           // mm_interconnect_0:onchip_d_memory_s2_write -> onchip_d_memory:write2
	wire  [31:0] mm_interconnect_0_onchip_d_memory_s2_writedata;                       // mm_interconnect_0:onchip_d_memory_s2_writedata -> onchip_d_memory:writedata2
	wire         mm_interconnect_0_onchip_d_memory_s2_clken;                           // mm_interconnect_0:onchip_d_memory_s2_clken -> onchip_d_memory:clken2
	wire  [31:0] nios2_gen2_0_data_master_readdata;                                    // mm_interconnect_1:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                                 // mm_interconnect_1:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                                 // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_1:nios2_gen2_0_data_master_debugaccess
	wire  [14:0] nios2_gen2_0_data_master_address;                                     // nios2_gen2_0:d_address -> mm_interconnect_1:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                                  // nios2_gen2_0:d_byteenable -> mm_interconnect_1:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                                        // nios2_gen2_0:d_read -> mm_interconnect_1:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_write;                                       // nios2_gen2_0:d_write -> mm_interconnect_1:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                                   // nios2_gen2_0:d_writedata -> mm_interconnect_1:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                             // mm_interconnect_1:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                          // mm_interconnect_1:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [14:0] nios2_gen2_0_instruction_master_address;                              // nios2_gen2_0:i_address -> mm_interconnect_1:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                                 // nios2_gen2_0:i_read -> mm_interconnect_1:nios2_gen2_0_instruction_master_read
	wire         mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_chipselect;           // mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_readdata;             // jtag_uart_0:av_readdata -> mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_waitrequest;          // jtag_uart_0:av_waitrequest -> mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_address;              // mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read;                 // mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write;                // mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_writedata;            // mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire         mm_interconnect_1_cnn_accelerator_avalon_0_avalon_slave_0_chipselect; // mm_interconnect_1:cnn_accelerator_avalon_0_avalon_slave_0_chipselect -> cnn_accelerator_avalon_0:AVS_s0_chipselect
	wire  [31:0] mm_interconnect_1_cnn_accelerator_avalon_0_avalon_slave_0_readdata;   // cnn_accelerator_avalon_0:AVS_s0_readdata -> mm_interconnect_1:cnn_accelerator_avalon_0_avalon_slave_0_readdata
	wire   [3:0] mm_interconnect_1_cnn_accelerator_avalon_0_avalon_slave_0_address;    // mm_interconnect_1:cnn_accelerator_avalon_0_avalon_slave_0_address -> cnn_accelerator_avalon_0:AVS_s0_adress
	wire         mm_interconnect_1_cnn_accelerator_avalon_0_avalon_slave_0_read;       // mm_interconnect_1:cnn_accelerator_avalon_0_avalon_slave_0_read -> cnn_accelerator_avalon_0:AVS_s0_read
	wire         mm_interconnect_1_cnn_accelerator_avalon_0_avalon_slave_0_write;      // mm_interconnect_1:cnn_accelerator_avalon_0_avalon_slave_0_write -> cnn_accelerator_avalon_0:AVS_s0_write
	wire  [31:0] mm_interconnect_1_cnn_accelerator_avalon_0_avalon_slave_0_writedata;  // mm_interconnect_1:cnn_accelerator_avalon_0_avalon_slave_0_writedata -> cnn_accelerator_avalon_0:AVS_s0_writedata
	wire  [31:0] mm_interconnect_1_nios2_gen2_0_debug_mem_slave_readdata;              // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_1:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_1_nios2_gen2_0_debug_mem_slave_waitrequest;           // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_1:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_1_nios2_gen2_0_debug_mem_slave_debugaccess;           // mm_interconnect_1:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_1_nios2_gen2_0_debug_mem_slave_address;               // mm_interconnect_1:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_1_nios2_gen2_0_debug_mem_slave_read;                  // mm_interconnect_1:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_1_nios2_gen2_0_debug_mem_slave_byteenable;            // mm_interconnect_1:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_1_nios2_gen2_0_debug_mem_slave_write;                 // mm_interconnect_1:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_1_nios2_gen2_0_debug_mem_slave_writedata;             // mm_interconnect_1:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire         mm_interconnect_1_onchip_ir_memory_s1_chipselect;                     // mm_interconnect_1:onchip_Ir_memory_s1_chipselect -> onchip_Ir_memory:chipselect
	wire  [31:0] mm_interconnect_1_onchip_ir_memory_s1_readdata;                       // onchip_Ir_memory:readdata -> mm_interconnect_1:onchip_Ir_memory_s1_readdata
	wire   [9:0] mm_interconnect_1_onchip_ir_memory_s1_address;                        // mm_interconnect_1:onchip_Ir_memory_s1_address -> onchip_Ir_memory:address
	wire   [3:0] mm_interconnect_1_onchip_ir_memory_s1_byteenable;                     // mm_interconnect_1:onchip_Ir_memory_s1_byteenable -> onchip_Ir_memory:byteenable
	wire         mm_interconnect_1_onchip_ir_memory_s1_write;                          // mm_interconnect_1:onchip_Ir_memory_s1_write -> onchip_Ir_memory:write
	wire  [31:0] mm_interconnect_1_onchip_ir_memory_s1_writedata;                      // mm_interconnect_1:onchip_Ir_memory_s1_writedata -> onchip_Ir_memory:writedata
	wire         mm_interconnect_1_onchip_ir_memory_s1_clken;                          // mm_interconnect_1:onchip_Ir_memory_s1_clken -> onchip_Ir_memory:clken
	wire         mm_interconnect_1_onchip_d_memory_s1_chipselect;                      // mm_interconnect_1:onchip_d_memory_s1_chipselect -> onchip_d_memory:chipselect
	wire  [31:0] mm_interconnect_1_onchip_d_memory_s1_readdata;                        // onchip_d_memory:readdata -> mm_interconnect_1:onchip_d_memory_s1_readdata
	wire   [9:0] mm_interconnect_1_onchip_d_memory_s1_address;                         // mm_interconnect_1:onchip_d_memory_s1_address -> onchip_d_memory:address
	wire   [3:0] mm_interconnect_1_onchip_d_memory_s1_byteenable;                      // mm_interconnect_1:onchip_d_memory_s1_byteenable -> onchip_d_memory:byteenable
	wire         mm_interconnect_1_onchip_d_memory_s1_write;                           // mm_interconnect_1:onchip_d_memory_s1_write -> onchip_d_memory:write
	wire  [31:0] mm_interconnect_1_onchip_d_memory_s1_writedata;                       // mm_interconnect_1:onchip_d_memory_s1_writedata -> onchip_d_memory:writedata
	wire         mm_interconnect_1_onchip_d_memory_s1_clken;                           // mm_interconnect_1:onchip_d_memory_s1_clken -> onchip_d_memory:clken
	wire         irq_mapper_receiver0_irq;                                             // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                                 // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                                       // rst_controller:reset_out -> [cnn_accelerator_avalon_0:AVS_Reset, jtag_uart_0:rst_n, mm_interconnect_0:cnn_accelerator_avalon_0_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_1:jtag_uart_0_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset;                                   // rst_controller_001:reset_out -> [irq_mapper:reset, mm_interconnect_0:onchip_d_memory_reset2_reset_bridge_in_reset_reset, mm_interconnect_1:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, onchip_Ir_memory:reset, onchip_d_memory:reset, onchip_d_memory:reset2, rst_translator:in_reset]
	wire         rst_controller_001_reset_out_reset_req;                               // rst_controller_001:reset_req -> [onchip_Ir_memory:reset_req, onchip_d_memory:reset_req, onchip_d_memory:reset_req2, rst_translator:reset_req_in]
	wire         nios2_gen2_0_debug_reset_request_reset;                               // nios2_gen2_0:debug_reset_request -> rst_controller_001:reset_in1

	ACCELERATOR_AVALON_INTERFACE #(
		.OFFMEM_DATA_WIDTH    (16),
		.OFFMEM_ADDR_WIDTH    (32),
		.BITWIDTH_DATA_OUT    (16),
		.BITWIDTH_IF_ROWS     (10),
		.BITWIDTH_IF_COLUMS   (11),
		.BITWIDTH_W_ROWS      (4),
		.BITWIDTH_W_COLUMS    (4),
		.BITWIDTH_IF_CHANNELS (2),
		.BITWIDTH_STRIDE      (4)
	) cnn_accelerator_avalon_0 (
		.AVS_s0_chipselect        (mm_interconnect_1_cnn_accelerator_avalon_0_avalon_slave_0_chipselect), //  avalon_slave_0.chipselect
		.AVS_s0_read              (mm_interconnect_1_cnn_accelerator_avalon_0_avalon_slave_0_read),       //                .read
		.AVS_s0_readdata          (mm_interconnect_1_cnn_accelerator_avalon_0_avalon_slave_0_readdata),   //                .readdata
		.AVS_s0_write             (mm_interconnect_1_cnn_accelerator_avalon_0_avalon_slave_0_write),      //                .write
		.AVS_s0_writedata         (mm_interconnect_1_cnn_accelerator_avalon_0_avalon_slave_0_writedata),  //                .writedata
		.AVS_s0_adress            (mm_interconnect_1_cnn_accelerator_avalon_0_avalon_slave_0_address),    //                .address
		.AVS_m0_adress            (cnn_accelerator_avalon_0_avalon_master_address),                       //   avalon_master.address
		.AVS_m0_byteenable        (cnn_accelerator_avalon_0_avalon_master_byteenable),                    //                .byteenable
		.AVS_m0_read              (cnn_accelerator_avalon_0_avalon_master_read),                          //                .read
		.AVS_m0_readdata          (cnn_accelerator_avalon_0_avalon_master_readdata),                      //                .readdata
		.AVS_m0_waitrequest       (cnn_accelerator_avalon_0_avalon_master_waitrequest),                   //                .waitrequest
		.AVS_m0_write             (cnn_accelerator_avalon_0_avalon_master_write),                         //                .write
		.AVS_m0_writedata         (cnn_accelerator_avalon_0_avalon_master_writedata),                     //                .writedata
		.AVS_Clk                  (clk_clk),                                                              //      clock_sink.clk
		.AVS_Reset                (~rst_controller_reset_out_reset),                                      //      reset_sink.reset_n
		.AVS_Counduit_Finished    (cnn_accelerator_avalon_0_control_signals_finished),                    // control_signals.finished
		.AVS_Counduit_Finished_Ok (cnn_accelerator_avalon_0_control_signals_finished_ok),                 //                .finished_ok
		.AVS_Counduit_Same_W      (cnn_accelerator_avalon_0_control_signals_same_w),                      //                .same_w
		.AVS_Counduit_Start       (cnn_accelerator_avalon_0_control_signals_start)                        //                .start
	);

	nios_system_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	nios_system_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                        //                     reset.reset_n
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	nios_system_onchip_Ir_memory onchip_ir_memory (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_1_onchip_ir_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_1_onchip_ir_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_1_onchip_ir_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_1_onchip_ir_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_1_onchip_ir_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_1_onchip_ir_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_1_onchip_ir_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),               // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req),           //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	nios_system_onchip_d_memory onchip_d_memory (
		.clk         (clk_clk),                                         //   clk1.clk
		.address     (mm_interconnect_1_onchip_d_memory_s1_address),    //     s1.address
		.clken       (mm_interconnect_1_onchip_d_memory_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_1_onchip_d_memory_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_1_onchip_d_memory_s1_write),      //       .write
		.readdata    (mm_interconnect_1_onchip_d_memory_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_1_onchip_d_memory_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_1_onchip_d_memory_s1_byteenable), //       .byteenable
		.reset       (rst_controller_001_reset_out_reset),              // reset1.reset
		.reset_req   (rst_controller_001_reset_out_reset_req),          //       .reset_req
		.address2    (mm_interconnect_0_onchip_d_memory_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_onchip_d_memory_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_onchip_d_memory_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_onchip_d_memory_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_onchip_d_memory_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_onchip_d_memory_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_onchip_d_memory_s2_byteenable), //       .byteenable
		.clk2        (clk_clk),                                         //   clk2.clk
		.reset2      (rst_controller_001_reset_out_reset),              // reset2.reset
		.reset_req2  (rst_controller_001_reset_out_reset_req),          //       .reset_req
		.freeze      (1'b0)                                             // (terminated)
	);

	nios_system_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                                   (clk_clk),                                            //                                                 clk_0_clk.clk
		.cnn_accelerator_avalon_0_reset_sink_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                     // cnn_accelerator_avalon_0_reset_sink_reset_bridge_in_reset.reset
		.onchip_d_memory_reset2_reset_bridge_in_reset_reset              (rst_controller_001_reset_out_reset),                 //              onchip_d_memory_reset2_reset_bridge_in_reset.reset
		.cnn_accelerator_avalon_0_avalon_master_address                  (cnn_accelerator_avalon_0_avalon_master_address),     //                    cnn_accelerator_avalon_0_avalon_master.address
		.cnn_accelerator_avalon_0_avalon_master_waitrequest              (cnn_accelerator_avalon_0_avalon_master_waitrequest), //                                                          .waitrequest
		.cnn_accelerator_avalon_0_avalon_master_byteenable               (cnn_accelerator_avalon_0_avalon_master_byteenable),  //                                                          .byteenable
		.cnn_accelerator_avalon_0_avalon_master_read                     (cnn_accelerator_avalon_0_avalon_master_read),        //                                                          .read
		.cnn_accelerator_avalon_0_avalon_master_readdata                 (cnn_accelerator_avalon_0_avalon_master_readdata),    //                                                          .readdata
		.cnn_accelerator_avalon_0_avalon_master_write                    (cnn_accelerator_avalon_0_avalon_master_write),       //                                                          .write
		.cnn_accelerator_avalon_0_avalon_master_writedata                (cnn_accelerator_avalon_0_avalon_master_writedata),   //                                                          .writedata
		.onchip_d_memory_s2_address                                      (mm_interconnect_0_onchip_d_memory_s2_address),       //                                        onchip_d_memory_s2.address
		.onchip_d_memory_s2_write                                        (mm_interconnect_0_onchip_d_memory_s2_write),         //                                                          .write
		.onchip_d_memory_s2_readdata                                     (mm_interconnect_0_onchip_d_memory_s2_readdata),      //                                                          .readdata
		.onchip_d_memory_s2_writedata                                    (mm_interconnect_0_onchip_d_memory_s2_writedata),     //                                                          .writedata
		.onchip_d_memory_s2_byteenable                                   (mm_interconnect_0_onchip_d_memory_s2_byteenable),    //                                                          .byteenable
		.onchip_d_memory_s2_chipselect                                   (mm_interconnect_0_onchip_d_memory_s2_chipselect),    //                                                          .chipselect
		.onchip_d_memory_s2_clken                                        (mm_interconnect_0_onchip_d_memory_s2_clken)          //                                                          .clken
	);

	nios_system_mm_interconnect_1 mm_interconnect_1 (
		.clk_0_clk_clk                                      (clk_clk),                                                              //                                clk_0_clk.clk
		.jtag_uart_0_reset_reset_bridge_in_reset_reset      (rst_controller_reset_out_reset),                                       //  jtag_uart_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset     (rst_controller_001_reset_out_reset),                                   // nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address                   (nios2_gen2_0_data_master_address),                                     //                 nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest               (nios2_gen2_0_data_master_waitrequest),                                 //                                         .waitrequest
		.nios2_gen2_0_data_master_byteenable                (nios2_gen2_0_data_master_byteenable),                                  //                                         .byteenable
		.nios2_gen2_0_data_master_read                      (nios2_gen2_0_data_master_read),                                        //                                         .read
		.nios2_gen2_0_data_master_readdata                  (nios2_gen2_0_data_master_readdata),                                    //                                         .readdata
		.nios2_gen2_0_data_master_write                     (nios2_gen2_0_data_master_write),                                       //                                         .write
		.nios2_gen2_0_data_master_writedata                 (nios2_gen2_0_data_master_writedata),                                   //                                         .writedata
		.nios2_gen2_0_data_master_debugaccess               (nios2_gen2_0_data_master_debugaccess),                                 //                                         .debugaccess
		.nios2_gen2_0_instruction_master_address            (nios2_gen2_0_instruction_master_address),                              //          nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest        (nios2_gen2_0_instruction_master_waitrequest),                          //                                         .waitrequest
		.nios2_gen2_0_instruction_master_read               (nios2_gen2_0_instruction_master_read),                                 //                                         .read
		.nios2_gen2_0_instruction_master_readdata           (nios2_gen2_0_instruction_master_readdata),                             //                                         .readdata
		.cnn_accelerator_avalon_0_avalon_slave_0_address    (mm_interconnect_1_cnn_accelerator_avalon_0_avalon_slave_0_address),    //  cnn_accelerator_avalon_0_avalon_slave_0.address
		.cnn_accelerator_avalon_0_avalon_slave_0_write      (mm_interconnect_1_cnn_accelerator_avalon_0_avalon_slave_0_write),      //                                         .write
		.cnn_accelerator_avalon_0_avalon_slave_0_read       (mm_interconnect_1_cnn_accelerator_avalon_0_avalon_slave_0_read),       //                                         .read
		.cnn_accelerator_avalon_0_avalon_slave_0_readdata   (mm_interconnect_1_cnn_accelerator_avalon_0_avalon_slave_0_readdata),   //                                         .readdata
		.cnn_accelerator_avalon_0_avalon_slave_0_writedata  (mm_interconnect_1_cnn_accelerator_avalon_0_avalon_slave_0_writedata),  //                                         .writedata
		.cnn_accelerator_avalon_0_avalon_slave_0_chipselect (mm_interconnect_1_cnn_accelerator_avalon_0_avalon_slave_0_chipselect), //                                         .chipselect
		.jtag_uart_0_avalon_jtag_slave_address              (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_address),              //            jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write                (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write),                //                                         .write
		.jtag_uart_0_avalon_jtag_slave_read                 (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read),                 //                                         .read
		.jtag_uart_0_avalon_jtag_slave_readdata             (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_readdata),             //                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata            (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_writedata),            //                                         .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest          (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_waitrequest),          //                                         .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect           (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_chipselect),           //                                         .chipselect
		.nios2_gen2_0_debug_mem_slave_address               (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_address),               //             nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write                 (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_write),                 //                                         .write
		.nios2_gen2_0_debug_mem_slave_read                  (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_read),                  //                                         .read
		.nios2_gen2_0_debug_mem_slave_readdata              (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_readdata),              //                                         .readdata
		.nios2_gen2_0_debug_mem_slave_writedata             (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_writedata),             //                                         .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable            (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_byteenable),            //                                         .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest           (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_waitrequest),           //                                         .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess           (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_debugaccess),           //                                         .debugaccess
		.onchip_d_memory_s1_address                         (mm_interconnect_1_onchip_d_memory_s1_address),                         //                       onchip_d_memory_s1.address
		.onchip_d_memory_s1_write                           (mm_interconnect_1_onchip_d_memory_s1_write),                           //                                         .write
		.onchip_d_memory_s1_readdata                        (mm_interconnect_1_onchip_d_memory_s1_readdata),                        //                                         .readdata
		.onchip_d_memory_s1_writedata                       (mm_interconnect_1_onchip_d_memory_s1_writedata),                       //                                         .writedata
		.onchip_d_memory_s1_byteenable                      (mm_interconnect_1_onchip_d_memory_s1_byteenable),                      //                                         .byteenable
		.onchip_d_memory_s1_chipselect                      (mm_interconnect_1_onchip_d_memory_s1_chipselect),                      //                                         .chipselect
		.onchip_d_memory_s1_clken                           (mm_interconnect_1_onchip_d_memory_s1_clken),                           //                                         .clken
		.onchip_Ir_memory_s1_address                        (mm_interconnect_1_onchip_ir_memory_s1_address),                        //                      onchip_Ir_memory_s1.address
		.onchip_Ir_memory_s1_write                          (mm_interconnect_1_onchip_ir_memory_s1_write),                          //                                         .write
		.onchip_Ir_memory_s1_readdata                       (mm_interconnect_1_onchip_ir_memory_s1_readdata),                       //                                         .readdata
		.onchip_Ir_memory_s1_writedata                      (mm_interconnect_1_onchip_ir_memory_s1_writedata),                      //                                         .writedata
		.onchip_Ir_memory_s1_byteenable                     (mm_interconnect_1_onchip_ir_memory_s1_byteenable),                     //                                         .byteenable
		.onchip_Ir_memory_s1_chipselect                     (mm_interconnect_1_onchip_ir_memory_s1_chipselect),                     //                                         .chipselect
		.onchip_Ir_memory_s1_clken                          (mm_interconnect_1_onchip_ir_memory_s1_clken)                           //                                         .clken
	);

	nios_system_irq_mapper irq_mapper (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.sender_irq    (nios2_gen2_0_irq_irq)                //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
