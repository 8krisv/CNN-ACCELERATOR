
module nios_system (
	clk_clk,
	cnn_accelerator_avalon_0_control_signals_finished,
	cnn_accelerator_avalon_0_control_signals_finished_ok,
	cnn_accelerator_avalon_0_control_signals_same_w,
	cnn_accelerator_avalon_0_control_signals_start,
	reset_reset_n);	

	input		clk_clk;
	output		cnn_accelerator_avalon_0_control_signals_finished;
	input		cnn_accelerator_avalon_0_control_signals_finished_ok;
	input		cnn_accelerator_avalon_0_control_signals_same_w;
	input		cnn_accelerator_avalon_0_control_signals_start;
	input		reset_reset_n;
endmodule
